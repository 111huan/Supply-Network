* layer: M1,VDD net: 0
R1 n1_0_0 n1_10_0 0.1
R2 n1_10_0 n1_20_0 0.1
R3 n1_0_10 n1_10_10 0.1
R4 n1_10_10 n1_20_10 0.1
R5 n1_0_20 n1_10_20 0.1
R6 n1_10_20 n1_20_20 0.1
* vias from: 0 to 3
V7 n1_0_0 n3_0_0 0.05
V8 n1_0_10 n3_0_10 0.05
V9 n1_0_20 n3_0_20 0.05
V10 n1_10_0 n3_10_0 0.05
V11 n1_10_10 n3_10_10 0.05
V12 n1_10_20 n3_10_20 0.05
V13 n1_20_0 n3_20_0 0.05
V14 n1_20_10 n3_20_10 0.05
V15 n1_20_20 n3_20_20 0.05
* layer: M2,VDD net: 3
R16 n3_0_0 n3_0_10 0.1
R17 n3_0_10 n3_0_20 0.1
R18 n3_10_0 n3_10_10 0.1
R19 n3_10_10 n3_10_20 0.1
R20 n3_20_0 n3_20_10 0.1
R21 n3_20_10 n3_20_20 0.1
rr22 n3_0_0 _X_n3_0_0 0
v22 _X_n3_0_0 0.5
rr23 n3_20_20 _X_n3_20_20 0
v23 _X_n3_20_20 0.5
iB0_0_v n1_0_0 0 0.03M
iB1_0_v n1_10_20 0 0.03M
