* layer: M1,VDD net: 0
R0 n0_0.0_0.0 n0_0.0001_0.0 0.014716220100000002
R1 n0_0.0001_0.0 n0_0.0002_0.0 0.014716220100000002
R2 n0_0.0002_0.0 n0_0.00030000000000000003_0.0 0.014716220100000002
R3 n0_0.00030000000000000003_0.0 n0_0.0004_0.0 0.014716220100000002
R4 n0_0.0004_0.0 n0_0.0005_0.0 0.014716220100000002
R5 n0_0.0005_0.0 n0_0.0006000000000000001_0.0 0.014716220100000002
R6 n0_0.0006000000000000001_0.0 n0_0.0007_0.0 0.014716220100000002
R7 n0_0.0007_0.0 n0_0.0008_0.0 0.014716220100000002
R8 n0_0.0008_0.0 n0_0.0009000000000000001_0.0 0.014716220100000002
R9 n0_0.0009000000000000001_0.0 n0_0.001_0.0 0.014716220100000002
R10 n0_0.001_0.0 n0_0.0011_0.0 0.014716220100000002
R11 n0_0.0011_0.0 n0_0.0012000000000000001_0.0 0.014716220100000002
R12 n0_0.0012000000000000001_0.0 n0_0.0013000000000000002_0.0 0.014716220100000002
R13 n0_0.0013000000000000002_0.0 n0_0.0014_0.0 0.014716220100000002
R14 n0_0.0014_0.0 n0_0.0015_0.0 0.014716220100000002
R15 n0_0.0015_0.0 n0_0.0016_0.0 0.014716220100000002
R16 n0_0.0_0.0001 n0_0.0001_0.0001 0.014716220100000002
R17 n0_0.0001_0.0001 n0_0.0002_0.0001 0.014716220100000002
R18 n0_0.0002_0.0001 n0_0.00030000000000000003_0.0001 0.014716220100000002
R19 n0_0.00030000000000000003_0.0001 n0_0.0004_0.0001 0.014716220100000002
R20 n0_0.0004_0.0001 n0_0.0005_0.0001 0.014716220100000002
R21 n0_0.0005_0.0001 n0_0.0006000000000000001_0.0001 0.014716220100000002
R22 n0_0.0006000000000000001_0.0001 n0_0.0007_0.0001 0.014716220100000002
R23 n0_0.0007_0.0001 n0_0.0008_0.0001 0.014716220100000002
R24 n0_0.0008_0.0001 n0_0.0009000000000000001_0.0001 0.014716220100000002
R25 n0_0.0009000000000000001_0.0001 n0_0.001_0.0001 0.014716220100000002
R26 n0_0.001_0.0001 n0_0.0011_0.0001 0.014716220100000002
R27 n0_0.0011_0.0001 n0_0.0012000000000000001_0.0001 0.014716220100000002
R28 n0_0.0012000000000000001_0.0001 n0_0.0013000000000000002_0.0001 0.014716220100000002
R29 n0_0.0013000000000000002_0.0001 n0_0.0014_0.0001 0.014716220100000002
R30 n0_0.0014_0.0001 n0_0.0015_0.0001 0.014716220100000002
R31 n0_0.0015_0.0001 n0_0.0016_0.0001 0.014716220100000002
R32 n0_0.0_0.0002 n0_0.0001_0.0002 0.014716220100000002
R33 n0_0.0001_0.0002 n0_0.0002_0.0002 0.014716220100000002
R34 n0_0.0002_0.0002 n0_0.00030000000000000003_0.0002 0.014716220100000002
R35 n0_0.00030000000000000003_0.0002 n0_0.0004_0.0002 0.014716220100000002
R36 n0_0.0004_0.0002 n0_0.0005_0.0002 0.014716220100000002
R37 n0_0.0005_0.0002 n0_0.0006000000000000001_0.0002 0.014716220100000002
R38 n0_0.0006000000000000001_0.0002 n0_0.0007_0.0002 0.014716220100000002
R39 n0_0.0007_0.0002 n0_0.0008_0.0002 0.014716220100000002
R40 n0_0.0008_0.0002 n0_0.0009000000000000001_0.0002 0.014716220100000002
R41 n0_0.0009000000000000001_0.0002 n0_0.001_0.0002 0.014716220100000002
R42 n0_0.001_0.0002 n0_0.0011_0.0002 0.014716220100000002
R43 n0_0.0011_0.0002 n0_0.0012000000000000001_0.0002 0.014716220100000002
R44 n0_0.0012000000000000001_0.0002 n0_0.0013000000000000002_0.0002 0.014716220100000002
R45 n0_0.0013000000000000002_0.0002 n0_0.0014_0.0002 0.014716220100000002
R46 n0_0.0014_0.0002 n0_0.0015_0.0002 0.014716220100000002
R47 n0_0.0015_0.0002 n0_0.0016_0.0002 0.014716220100000002
R48 n0_0.0_0.00030000000000000003 n0_0.0001_0.00030000000000000003 0.014716220100000002
R49 n0_0.0001_0.00030000000000000003 n0_0.0002_0.00030000000000000003 0.014716220100000002
R50 n0_0.0002_0.00030000000000000003 n0_0.00030000000000000003_0.00030000000000000003 0.014716220100000002
R51 n0_0.00030000000000000003_0.00030000000000000003 n0_0.0004_0.00030000000000000003 0.014716220100000002
R52 n0_0.0004_0.00030000000000000003 n0_0.0005_0.00030000000000000003 0.014716220100000002
R53 n0_0.0005_0.00030000000000000003 n0_0.0006000000000000001_0.00030000000000000003 0.014716220100000002
R54 n0_0.0006000000000000001_0.00030000000000000003 n0_0.0007_0.00030000000000000003 0.014716220100000002
R55 n0_0.0007_0.00030000000000000003 n0_0.0008_0.00030000000000000003 0.014716220100000002
R56 n0_0.0008_0.00030000000000000003 n0_0.0009000000000000001_0.00030000000000000003 0.014716220100000002
R57 n0_0.0009000000000000001_0.00030000000000000003 n0_0.001_0.00030000000000000003 0.014716220100000002
R58 n0_0.001_0.00030000000000000003 n0_0.0011_0.00030000000000000003 0.014716220100000002
R59 n0_0.0011_0.00030000000000000003 n0_0.0012000000000000001_0.00030000000000000003 0.014716220100000002
R60 n0_0.0012000000000000001_0.00030000000000000003 n0_0.0013000000000000002_0.00030000000000000003 0.014716220100000002
R61 n0_0.0013000000000000002_0.00030000000000000003 n0_0.0014_0.00030000000000000003 0.014716220100000002
R62 n0_0.0014_0.00030000000000000003 n0_0.0015_0.00030000000000000003 0.014716220100000002
R63 n0_0.0015_0.00030000000000000003 n0_0.0016_0.00030000000000000003 0.014716220100000002
R64 n0_0.0_0.0004 n0_0.0001_0.0004 0.014716220100000002
R65 n0_0.0001_0.0004 n0_0.0002_0.0004 0.014716220100000002
R66 n0_0.0002_0.0004 n0_0.00030000000000000003_0.0004 0.014716220100000002
R67 n0_0.00030000000000000003_0.0004 n0_0.0004_0.0004 0.014716220100000002
R68 n0_0.0004_0.0004 n0_0.0005_0.0004 0.014716220100000002
R69 n0_0.0005_0.0004 n0_0.0006000000000000001_0.0004 0.014716220100000002
R70 n0_0.0006000000000000001_0.0004 n0_0.0007_0.0004 0.014716220100000002
R71 n0_0.0007_0.0004 n0_0.0008_0.0004 0.014716220100000002
R72 n0_0.0008_0.0004 n0_0.0009000000000000001_0.0004 0.014716220100000002
R73 n0_0.0009000000000000001_0.0004 n0_0.001_0.0004 0.014716220100000002
R74 n0_0.001_0.0004 n0_0.0011_0.0004 0.014716220100000002
R75 n0_0.0011_0.0004 n0_0.0012000000000000001_0.0004 0.014716220100000002
R76 n0_0.0012000000000000001_0.0004 n0_0.0013000000000000002_0.0004 0.014716220100000002
R77 n0_0.0013000000000000002_0.0004 n0_0.0014_0.0004 0.014716220100000002
R78 n0_0.0014_0.0004 n0_0.0015_0.0004 0.014716220100000002
R79 n0_0.0015_0.0004 n0_0.0016_0.0004 0.014716220100000002
R80 n0_0.0_0.0005 n0_0.0001_0.0005 0.014716220100000002
R81 n0_0.0001_0.0005 n0_0.0002_0.0005 0.014716220100000002
R82 n0_0.0002_0.0005 n0_0.00030000000000000003_0.0005 0.014716220100000002
R83 n0_0.00030000000000000003_0.0005 n0_0.0004_0.0005 0.014716220100000002
R84 n0_0.0004_0.0005 n0_0.0005_0.0005 0.014716220100000002
R85 n0_0.0005_0.0005 n0_0.0006000000000000001_0.0005 0.014716220100000002
R86 n0_0.0006000000000000001_0.0005 n0_0.0007_0.0005 0.014716220100000002
R87 n0_0.0007_0.0005 n0_0.0008_0.0005 0.014716220100000002
R88 n0_0.0008_0.0005 n0_0.0009000000000000001_0.0005 0.014716220100000002
R89 n0_0.0009000000000000001_0.0005 n0_0.001_0.0005 0.014716220100000002
R90 n0_0.001_0.0005 n0_0.0011_0.0005 0.014716220100000002
R91 n0_0.0011_0.0005 n0_0.0012000000000000001_0.0005 0.014716220100000002
R92 n0_0.0012000000000000001_0.0005 n0_0.0013000000000000002_0.0005 0.014716220100000002
R93 n0_0.0013000000000000002_0.0005 n0_0.0014_0.0005 0.014716220100000002
R94 n0_0.0014_0.0005 n0_0.0015_0.0005 0.014716220100000002
R95 n0_0.0015_0.0005 n0_0.0016_0.0005 0.014716220100000002
R96 n0_0.0_0.0006000000000000001 n0_0.0001_0.0006000000000000001 0.014716220100000002
R97 n0_0.0001_0.0006000000000000001 n0_0.0002_0.0006000000000000001 0.014716220100000002
R98 n0_0.0002_0.0006000000000000001 n0_0.00030000000000000003_0.0006000000000000001 0.014716220100000002
R99 n0_0.00030000000000000003_0.0006000000000000001 n0_0.0004_0.0006000000000000001 0.014716220100000002
R100 n0_0.0004_0.0006000000000000001 n0_0.0005_0.0006000000000000001 0.014716220100000002
R101 n0_0.0005_0.0006000000000000001 n0_0.0006000000000000001_0.0006000000000000001 0.014716220100000002
R102 n0_0.0006000000000000001_0.0006000000000000001 n0_0.0007_0.0006000000000000001 0.014716220100000002
R103 n0_0.0007_0.0006000000000000001 n0_0.0008_0.0006000000000000001 0.014716220100000002
R104 n0_0.0008_0.0006000000000000001 n0_0.0009000000000000001_0.0006000000000000001 0.014716220100000002
R105 n0_0.0009000000000000001_0.0006000000000000001 n0_0.001_0.0006000000000000001 0.014716220100000002
R106 n0_0.001_0.0006000000000000001 n0_0.0011_0.0006000000000000001 0.014716220100000002
R107 n0_0.0011_0.0006000000000000001 n0_0.0012000000000000001_0.0006000000000000001 0.014716220100000002
R108 n0_0.0012000000000000001_0.0006000000000000001 n0_0.0013000000000000002_0.0006000000000000001 0.014716220100000002
R109 n0_0.0013000000000000002_0.0006000000000000001 n0_0.0014_0.0006000000000000001 0.014716220100000002
R110 n0_0.0014_0.0006000000000000001 n0_0.0015_0.0006000000000000001 0.014716220100000002
R111 n0_0.0015_0.0006000000000000001 n0_0.0016_0.0006000000000000001 0.014716220100000002
R112 n0_0.0_0.0007 n0_0.0001_0.0007 0.014716220100000002
R113 n0_0.0001_0.0007 n0_0.0002_0.0007 0.014716220100000002
R114 n0_0.0002_0.0007 n0_0.00030000000000000003_0.0007 0.014716220100000002
R115 n0_0.00030000000000000003_0.0007 n0_0.0004_0.0007 0.014716220100000002
R116 n0_0.0004_0.0007 n0_0.0005_0.0007 0.014716220100000002
R117 n0_0.0005_0.0007 n0_0.0006000000000000001_0.0007 0.014716220100000002
R118 n0_0.0006000000000000001_0.0007 n0_0.0007_0.0007 0.014716220100000002
R119 n0_0.0007_0.0007 n0_0.0008_0.0007 0.014716220100000002
R120 n0_0.0008_0.0007 n0_0.0009000000000000001_0.0007 0.014716220100000002
R121 n0_0.0009000000000000001_0.0007 n0_0.001_0.0007 0.014716220100000002
R122 n0_0.001_0.0007 n0_0.0011_0.0007 0.014716220100000002
R123 n0_0.0011_0.0007 n0_0.0012000000000000001_0.0007 0.014716220100000002
R124 n0_0.0012000000000000001_0.0007 n0_0.0013000000000000002_0.0007 0.014716220100000002
R125 n0_0.0013000000000000002_0.0007 n0_0.0014_0.0007 0.014716220100000002
R126 n0_0.0014_0.0007 n0_0.0015_0.0007 0.014716220100000002
R127 n0_0.0015_0.0007 n0_0.0016_0.0007 0.014716220100000002
R128 n0_0.0_0.0008 n0_0.0001_0.0008 0.014716220100000002
R129 n0_0.0001_0.0008 n0_0.0002_0.0008 0.014716220100000002
R130 n0_0.0002_0.0008 n0_0.00030000000000000003_0.0008 0.014716220100000002
R131 n0_0.00030000000000000003_0.0008 n0_0.0004_0.0008 0.014716220100000002
R132 n0_0.0004_0.0008 n0_0.0005_0.0008 0.014716220100000002
R133 n0_0.0005_0.0008 n0_0.0006000000000000001_0.0008 0.014716220100000002
R134 n0_0.0006000000000000001_0.0008 n0_0.0007_0.0008 0.014716220100000002
R135 n0_0.0007_0.0008 n0_0.0008_0.0008 0.014716220100000002
R136 n0_0.0008_0.0008 n0_0.0009000000000000001_0.0008 0.014716220100000002
R137 n0_0.0009000000000000001_0.0008 n0_0.001_0.0008 0.014716220100000002
R138 n0_0.001_0.0008 n0_0.0011_0.0008 0.014716220100000002
R139 n0_0.0011_0.0008 n0_0.0012000000000000001_0.0008 0.014716220100000002
R140 n0_0.0012000000000000001_0.0008 n0_0.0013000000000000002_0.0008 0.014716220100000002
R141 n0_0.0013000000000000002_0.0008 n0_0.0014_0.0008 0.014716220100000002
R142 n0_0.0014_0.0008 n0_0.0015_0.0008 0.014716220100000002
R143 n0_0.0015_0.0008 n0_0.0016_0.0008 0.014716220100000002
R144 n0_0.0_0.0009000000000000001 n0_0.0001_0.0009000000000000001 0.014716220100000002
R145 n0_0.0001_0.0009000000000000001 n0_0.0002_0.0009000000000000001 0.014716220100000002
R146 n0_0.0002_0.0009000000000000001 n0_0.00030000000000000003_0.0009000000000000001 0.014716220100000002
R147 n0_0.00030000000000000003_0.0009000000000000001 n0_0.0004_0.0009000000000000001 0.014716220100000002
R148 n0_0.0004_0.0009000000000000001 n0_0.0005_0.0009000000000000001 0.014716220100000002
R149 n0_0.0005_0.0009000000000000001 n0_0.0006000000000000001_0.0009000000000000001 0.014716220100000002
R150 n0_0.0006000000000000001_0.0009000000000000001 n0_0.0007_0.0009000000000000001 0.014716220100000002
R151 n0_0.0007_0.0009000000000000001 n0_0.0008_0.0009000000000000001 0.014716220100000002
R152 n0_0.0008_0.0009000000000000001 n0_0.0009000000000000001_0.0009000000000000001 0.014716220100000002
R153 n0_0.0009000000000000001_0.0009000000000000001 n0_0.001_0.0009000000000000001 0.014716220100000002
R154 n0_0.001_0.0009000000000000001 n0_0.0011_0.0009000000000000001 0.014716220100000002
R155 n0_0.0011_0.0009000000000000001 n0_0.0012000000000000001_0.0009000000000000001 0.014716220100000002
R156 n0_0.0012000000000000001_0.0009000000000000001 n0_0.0013000000000000002_0.0009000000000000001 0.014716220100000002
R157 n0_0.0013000000000000002_0.0009000000000000001 n0_0.0014_0.0009000000000000001 0.014716220100000002
R158 n0_0.0014_0.0009000000000000001 n0_0.0015_0.0009000000000000001 0.014716220100000002
R159 n0_0.0015_0.0009000000000000001 n0_0.0016_0.0009000000000000001 0.014716220100000002
R160 n0_0.0_0.001 n0_0.0001_0.001 0.014716220100000002
R161 n0_0.0001_0.001 n0_0.0002_0.001 0.014716220100000002
R162 n0_0.0002_0.001 n0_0.00030000000000000003_0.001 0.014716220100000002
R163 n0_0.00030000000000000003_0.001 n0_0.0004_0.001 0.014716220100000002
R164 n0_0.0004_0.001 n0_0.0005_0.001 0.014716220100000002
R165 n0_0.0005_0.001 n0_0.0006000000000000001_0.001 0.014716220100000002
R166 n0_0.0006000000000000001_0.001 n0_0.0007_0.001 0.014716220100000002
R167 n0_0.0007_0.001 n0_0.0008_0.001 0.014716220100000002
R168 n0_0.0008_0.001 n0_0.0009000000000000001_0.001 0.014716220100000002
R169 n0_0.0009000000000000001_0.001 n0_0.001_0.001 0.014716220100000002
R170 n0_0.001_0.001 n0_0.0011_0.001 0.014716220100000002
R171 n0_0.0011_0.001 n0_0.0012000000000000001_0.001 0.014716220100000002
R172 n0_0.0012000000000000001_0.001 n0_0.0013000000000000002_0.001 0.014716220100000002
R173 n0_0.0013000000000000002_0.001 n0_0.0014_0.001 0.014716220100000002
R174 n0_0.0014_0.001 n0_0.0015_0.001 0.014716220100000002
R175 n0_0.0015_0.001 n0_0.0016_0.001 0.014716220100000002
R176 n0_0.0_0.0011 n0_0.0001_0.0011 0.014716220100000002
R177 n0_0.0001_0.0011 n0_0.0002_0.0011 0.014716220100000002
R178 n0_0.0002_0.0011 n0_0.00030000000000000003_0.0011 0.014716220100000002
R179 n0_0.00030000000000000003_0.0011 n0_0.0004_0.0011 0.014716220100000002
R180 n0_0.0004_0.0011 n0_0.0005_0.0011 0.014716220100000002
R181 n0_0.0005_0.0011 n0_0.0006000000000000001_0.0011 0.014716220100000002
R182 n0_0.0006000000000000001_0.0011 n0_0.0007_0.0011 0.014716220100000002
R183 n0_0.0007_0.0011 n0_0.0008_0.0011 0.014716220100000002
R184 n0_0.0008_0.0011 n0_0.0009000000000000001_0.0011 0.014716220100000002
R185 n0_0.0009000000000000001_0.0011 n0_0.001_0.0011 0.014716220100000002
R186 n0_0.001_0.0011 n0_0.0011_0.0011 0.014716220100000002
R187 n0_0.0011_0.0011 n0_0.0012000000000000001_0.0011 0.014716220100000002
R188 n0_0.0012000000000000001_0.0011 n0_0.0013000000000000002_0.0011 0.014716220100000002
R189 n0_0.0013000000000000002_0.0011 n0_0.0014_0.0011 0.014716220100000002
R190 n0_0.0014_0.0011 n0_0.0015_0.0011 0.014716220100000002
R191 n0_0.0015_0.0011 n0_0.0016_0.0011 0.014716220100000002
R192 n0_0.0_0.0012000000000000001 n0_0.0001_0.0012000000000000001 0.014716220100000002
R193 n0_0.0001_0.0012000000000000001 n0_0.0002_0.0012000000000000001 0.014716220100000002
R194 n0_0.0002_0.0012000000000000001 n0_0.00030000000000000003_0.0012000000000000001 0.014716220100000002
R195 n0_0.00030000000000000003_0.0012000000000000001 n0_0.0004_0.0012000000000000001 0.014716220100000002
R196 n0_0.0004_0.0012000000000000001 n0_0.0005_0.0012000000000000001 0.014716220100000002
R197 n0_0.0005_0.0012000000000000001 n0_0.0006000000000000001_0.0012000000000000001 0.014716220100000002
R198 n0_0.0006000000000000001_0.0012000000000000001 n0_0.0007_0.0012000000000000001 0.014716220100000002
R199 n0_0.0007_0.0012000000000000001 n0_0.0008_0.0012000000000000001 0.014716220100000002
R200 n0_0.0008_0.0012000000000000001 n0_0.0009000000000000001_0.0012000000000000001 0.014716220100000002
R201 n0_0.0009000000000000001_0.0012000000000000001 n0_0.001_0.0012000000000000001 0.014716220100000002
R202 n0_0.001_0.0012000000000000001 n0_0.0011_0.0012000000000000001 0.014716220100000002
R203 n0_0.0011_0.0012000000000000001 n0_0.0012000000000000001_0.0012000000000000001 0.014716220100000002
R204 n0_0.0012000000000000001_0.0012000000000000001 n0_0.0013000000000000002_0.0012000000000000001 0.014716220100000002
R205 n0_0.0013000000000000002_0.0012000000000000001 n0_0.0014_0.0012000000000000001 0.014716220100000002
R206 n0_0.0014_0.0012000000000000001 n0_0.0015_0.0012000000000000001 0.014716220100000002
R207 n0_0.0015_0.0012000000000000001 n0_0.0016_0.0012000000000000001 0.014716220100000002
R208 n0_0.0_0.0013000000000000002 n0_0.0001_0.0013000000000000002 0.014716220100000002
R209 n0_0.0001_0.0013000000000000002 n0_0.0002_0.0013000000000000002 0.014716220100000002
R210 n0_0.0002_0.0013000000000000002 n0_0.00030000000000000003_0.0013000000000000002 0.014716220100000002
R211 n0_0.00030000000000000003_0.0013000000000000002 n0_0.0004_0.0013000000000000002 0.014716220100000002
R212 n0_0.0004_0.0013000000000000002 n0_0.0005_0.0013000000000000002 0.014716220100000002
R213 n0_0.0005_0.0013000000000000002 n0_0.0006000000000000001_0.0013000000000000002 0.014716220100000002
R214 n0_0.0006000000000000001_0.0013000000000000002 n0_0.0007_0.0013000000000000002 0.014716220100000002
R215 n0_0.0007_0.0013000000000000002 n0_0.0008_0.0013000000000000002 0.014716220100000002
R216 n0_0.0008_0.0013000000000000002 n0_0.0009000000000000001_0.0013000000000000002 0.014716220100000002
R217 n0_0.0009000000000000001_0.0013000000000000002 n0_0.001_0.0013000000000000002 0.014716220100000002
R218 n0_0.001_0.0013000000000000002 n0_0.0011_0.0013000000000000002 0.014716220100000002
R219 n0_0.0011_0.0013000000000000002 n0_0.0012000000000000001_0.0013000000000000002 0.014716220100000002
R220 n0_0.0012000000000000001_0.0013000000000000002 n0_0.0013000000000000002_0.0013000000000000002 0.014716220100000002
R221 n0_0.0013000000000000002_0.0013000000000000002 n0_0.0014_0.0013000000000000002 0.014716220100000002
R222 n0_0.0014_0.0013000000000000002 n0_0.0015_0.0013000000000000002 0.014716220100000002
R223 n0_0.0015_0.0013000000000000002 n0_0.0016_0.0013000000000000002 0.014716220100000002
R224 n0_0.0_0.0014 n0_0.0001_0.0014 0.014716220100000002
R225 n0_0.0001_0.0014 n0_0.0002_0.0014 0.014716220100000002
R226 n0_0.0002_0.0014 n0_0.00030000000000000003_0.0014 0.014716220100000002
R227 n0_0.00030000000000000003_0.0014 n0_0.0004_0.0014 0.014716220100000002
R228 n0_0.0004_0.0014 n0_0.0005_0.0014 0.014716220100000002
R229 n0_0.0005_0.0014 n0_0.0006000000000000001_0.0014 0.014716220100000002
R230 n0_0.0006000000000000001_0.0014 n0_0.0007_0.0014 0.014716220100000002
R231 n0_0.0007_0.0014 n0_0.0008_0.0014 0.014716220100000002
R232 n0_0.0008_0.0014 n0_0.0009000000000000001_0.0014 0.014716220100000002
R233 n0_0.0009000000000000001_0.0014 n0_0.001_0.0014 0.014716220100000002
R234 n0_0.001_0.0014 n0_0.0011_0.0014 0.014716220100000002
R235 n0_0.0011_0.0014 n0_0.0012000000000000001_0.0014 0.014716220100000002
R236 n0_0.0012000000000000001_0.0014 n0_0.0013000000000000002_0.0014 0.014716220100000002
R237 n0_0.0013000000000000002_0.0014 n0_0.0014_0.0014 0.014716220100000002
R238 n0_0.0014_0.0014 n0_0.0015_0.0014 0.014716220100000002
R239 n0_0.0015_0.0014 n0_0.0016_0.0014 0.014716220100000002
R240 n0_0.0_0.0015 n0_0.0001_0.0015 0.014716220100000002
R241 n0_0.0001_0.0015 n0_0.0002_0.0015 0.014716220100000002
R242 n0_0.0002_0.0015 n0_0.00030000000000000003_0.0015 0.014716220100000002
R243 n0_0.00030000000000000003_0.0015 n0_0.0004_0.0015 0.014716220100000002
R244 n0_0.0004_0.0015 n0_0.0005_0.0015 0.014716220100000002
R245 n0_0.0005_0.0015 n0_0.0006000000000000001_0.0015 0.014716220100000002
R246 n0_0.0006000000000000001_0.0015 n0_0.0007_0.0015 0.014716220100000002
R247 n0_0.0007_0.0015 n0_0.0008_0.0015 0.014716220100000002
R248 n0_0.0008_0.0015 n0_0.0009000000000000001_0.0015 0.014716220100000002
R249 n0_0.0009000000000000001_0.0015 n0_0.001_0.0015 0.014716220100000002
R250 n0_0.001_0.0015 n0_0.0011_0.0015 0.014716220100000002
R251 n0_0.0011_0.0015 n0_0.0012000000000000001_0.0015 0.014716220100000002
R252 n0_0.0012000000000000001_0.0015 n0_0.0013000000000000002_0.0015 0.014716220100000002
R253 n0_0.0013000000000000002_0.0015 n0_0.0014_0.0015 0.014716220100000002
R254 n0_0.0014_0.0015 n0_0.0015_0.0015 0.014716220100000002
R255 n0_0.0015_0.0015 n0_0.0016_0.0015 0.014716220100000002
R256 n0_0.0_0.0016 n0_0.0001_0.0016 0.014716220100000002
R257 n0_0.0001_0.0016 n0_0.0002_0.0016 0.014716220100000002
R258 n0_0.0002_0.0016 n0_0.00030000000000000003_0.0016 0.014716220100000002
R259 n0_0.00030000000000000003_0.0016 n0_0.0004_0.0016 0.014716220100000002
R260 n0_0.0004_0.0016 n0_0.0005_0.0016 0.014716220100000002
R261 n0_0.0005_0.0016 n0_0.0006000000000000001_0.0016 0.014716220100000002
R262 n0_0.0006000000000000001_0.0016 n0_0.0007_0.0016 0.014716220100000002
R263 n0_0.0007_0.0016 n0_0.0008_0.0016 0.014716220100000002
R264 n0_0.0008_0.0016 n0_0.0009000000000000001_0.0016 0.014716220100000002
R265 n0_0.0009000000000000001_0.0016 n0_0.001_0.0016 0.014716220100000002
R266 n0_0.001_0.0016 n0_0.0011_0.0016 0.014716220100000002
R267 n0_0.0011_0.0016 n0_0.0012000000000000001_0.0016 0.014716220100000002
R268 n0_0.0012000000000000001_0.0016 n0_0.0013000000000000002_0.0016 0.014716220100000002
R269 n0_0.0013000000000000002_0.0016 n0_0.0014_0.0016 0.014716220100000002
R270 n0_0.0014_0.0016 n0_0.0015_0.0016 0.014716220100000002
R271 n0_0.0015_0.0016 n0_0.0016_0.0016 0.014716220100000002
* vias from: 0 to 2
V272 n0_0.0_0.0 n2_0.0_0.0 0
V273 n0_0.0_0.0001 n2_0.0_0.0001 0
V274 n0_0.0_0.0002 n2_0.0_0.0002 0
V275 n0_0.0_0.00030000000000000003 n2_0.0_0.00030000000000000003 0
V276 n0_0.0_0.0004 n2_0.0_0.0004 0
V277 n0_0.0_0.0005 n2_0.0_0.0005 0
V278 n0_0.0_0.0006000000000000001 n2_0.0_0.0006000000000000001 0
V279 n0_0.0_0.0007 n2_0.0_0.0007 0
V280 n0_0.0_0.0008 n2_0.0_0.0008 0
V281 n0_0.0_0.0009000000000000001 n2_0.0_0.0009000000000000001 0
V282 n0_0.0_0.001 n2_0.0_0.001 0
V283 n0_0.0_0.0011 n2_0.0_0.0011 0
V284 n0_0.0_0.0012000000000000001 n2_0.0_0.0012000000000000001 0
V285 n0_0.0_0.0013000000000000002 n2_0.0_0.0013000000000000002 0
V286 n0_0.0_0.0014 n2_0.0_0.0014 0
V287 n0_0.0_0.0015 n2_0.0_0.0015 0
V288 n0_0.0_0.0016 n2_0.0_0.0016 0
V289 n0_0.0002_0.0 n2_0.0002_0.0 0
V290 n0_0.0002_0.0001 n2_0.0002_0.0001 0
V291 n0_0.0002_0.0002 n2_0.0002_0.0002 0
V292 n0_0.0002_0.00030000000000000003 n2_0.0002_0.00030000000000000003 0
V293 n0_0.0002_0.0004 n2_0.0002_0.0004 0
V294 n0_0.0002_0.0005 n2_0.0002_0.0005 0
V295 n0_0.0002_0.0006000000000000001 n2_0.0002_0.0006000000000000001 0
V296 n0_0.0002_0.0007 n2_0.0002_0.0007 0
V297 n0_0.0002_0.0008 n2_0.0002_0.0008 0
V298 n0_0.0002_0.0009000000000000001 n2_0.0002_0.0009000000000000001 0
V299 n0_0.0002_0.001 n2_0.0002_0.001 0
V300 n0_0.0002_0.0011 n2_0.0002_0.0011 0
V301 n0_0.0002_0.0012000000000000001 n2_0.0002_0.0012000000000000001 0
V302 n0_0.0002_0.0013000000000000002 n2_0.0002_0.0013000000000000002 0
V303 n0_0.0002_0.0014 n2_0.0002_0.0014 0
V304 n0_0.0002_0.0015 n2_0.0002_0.0015 0
V305 n0_0.0002_0.0016 n2_0.0002_0.0016 0
V306 n0_0.0004_0.0 n2_0.0004_0.0 0
V307 n0_0.0004_0.0001 n2_0.0004_0.0001 0
V308 n0_0.0004_0.0002 n2_0.0004_0.0002 0
V309 n0_0.0004_0.00030000000000000003 n2_0.0004_0.00030000000000000003 0
V310 n0_0.0004_0.0004 n2_0.0004_0.0004 0
V311 n0_0.0004_0.0005 n2_0.0004_0.0005 0
V312 n0_0.0004_0.0006000000000000001 n2_0.0004_0.0006000000000000001 0
V313 n0_0.0004_0.0007 n2_0.0004_0.0007 0
V314 n0_0.0004_0.0008 n2_0.0004_0.0008 0
V315 n0_0.0004_0.0009000000000000001 n2_0.0004_0.0009000000000000001 0
V316 n0_0.0004_0.001 n2_0.0004_0.001 0
V317 n0_0.0004_0.0011 n2_0.0004_0.0011 0
V318 n0_0.0004_0.0012000000000000001 n2_0.0004_0.0012000000000000001 0
V319 n0_0.0004_0.0013000000000000002 n2_0.0004_0.0013000000000000002 0
V320 n0_0.0004_0.0014 n2_0.0004_0.0014 0
V321 n0_0.0004_0.0015 n2_0.0004_0.0015 0
V322 n0_0.0004_0.0016 n2_0.0004_0.0016 0
V323 n0_0.0006000000000000001_0.0 n2_0.0006000000000000001_0.0 0
V324 n0_0.0006000000000000001_0.0001 n2_0.0006000000000000001_0.0001 0
V325 n0_0.0006000000000000001_0.0002 n2_0.0006000000000000001_0.0002 0
V326 n0_0.0006000000000000001_0.00030000000000000003 n2_0.0006000000000000001_0.00030000000000000003 0
V327 n0_0.0006000000000000001_0.0004 n2_0.0006000000000000001_0.0004 0
V328 n0_0.0006000000000000001_0.0005 n2_0.0006000000000000001_0.0005 0
V329 n0_0.0006000000000000001_0.0006000000000000001 n2_0.0006000000000000001_0.0006000000000000001 0
V330 n0_0.0006000000000000001_0.0007 n2_0.0006000000000000001_0.0007 0
V331 n0_0.0006000000000000001_0.0008 n2_0.0006000000000000001_0.0008 0
V332 n0_0.0006000000000000001_0.0009000000000000001 n2_0.0006000000000000001_0.0009000000000000001 0
V333 n0_0.0006000000000000001_0.001 n2_0.0006000000000000001_0.001 0
V334 n0_0.0006000000000000001_0.0011 n2_0.0006000000000000001_0.0011 0
V335 n0_0.0006000000000000001_0.0012000000000000001 n2_0.0006000000000000001_0.0012000000000000001 0
V336 n0_0.0006000000000000001_0.0013000000000000002 n2_0.0006000000000000001_0.0013000000000000002 0
V337 n0_0.0006000000000000001_0.0014 n2_0.0006000000000000001_0.0014 0
V338 n0_0.0006000000000000001_0.0015 n2_0.0006000000000000001_0.0015 0
V339 n0_0.0006000000000000001_0.0016 n2_0.0006000000000000001_0.0016 0
V340 n0_0.0008_0.0 n2_0.0008_0.0 0
V341 n0_0.0008_0.0001 n2_0.0008_0.0001 0
V342 n0_0.0008_0.0002 n2_0.0008_0.0002 0
V343 n0_0.0008_0.00030000000000000003 n2_0.0008_0.00030000000000000003 0
V344 n0_0.0008_0.0004 n2_0.0008_0.0004 0
V345 n0_0.0008_0.0005 n2_0.0008_0.0005 0
V346 n0_0.0008_0.0006000000000000001 n2_0.0008_0.0006000000000000001 0
V347 n0_0.0008_0.0007 n2_0.0008_0.0007 0
V348 n0_0.0008_0.0008 n2_0.0008_0.0008 0
V349 n0_0.0008_0.0009000000000000001 n2_0.0008_0.0009000000000000001 0
V350 n0_0.0008_0.001 n2_0.0008_0.001 0
V351 n0_0.0008_0.0011 n2_0.0008_0.0011 0
V352 n0_0.0008_0.0012000000000000001 n2_0.0008_0.0012000000000000001 0
V353 n0_0.0008_0.0013000000000000002 n2_0.0008_0.0013000000000000002 0
V354 n0_0.0008_0.0014 n2_0.0008_0.0014 0
V355 n0_0.0008_0.0015 n2_0.0008_0.0015 0
V356 n0_0.0008_0.0016 n2_0.0008_0.0016 0
V357 n0_0.001_0.0 n2_0.001_0.0 0
V358 n0_0.001_0.0001 n2_0.001_0.0001 0
V359 n0_0.001_0.0002 n2_0.001_0.0002 0
V360 n0_0.001_0.00030000000000000003 n2_0.001_0.00030000000000000003 0
V361 n0_0.001_0.0004 n2_0.001_0.0004 0
V362 n0_0.001_0.0005 n2_0.001_0.0005 0
V363 n0_0.001_0.0006000000000000001 n2_0.001_0.0006000000000000001 0
V364 n0_0.001_0.0007 n2_0.001_0.0007 0
V365 n0_0.001_0.0008 n2_0.001_0.0008 0
V366 n0_0.001_0.0009000000000000001 n2_0.001_0.0009000000000000001 0
V367 n0_0.001_0.001 n2_0.001_0.001 0
V368 n0_0.001_0.0011 n2_0.001_0.0011 0
V369 n0_0.001_0.0012000000000000001 n2_0.001_0.0012000000000000001 0
V370 n0_0.001_0.0013000000000000002 n2_0.001_0.0013000000000000002 0
V371 n0_0.001_0.0014 n2_0.001_0.0014 0
V372 n0_0.001_0.0015 n2_0.001_0.0015 0
V373 n0_0.001_0.0016 n2_0.001_0.0016 0
V374 n0_0.0012000000000000001_0.0 n2_0.0012000000000000001_0.0 0
V375 n0_0.0012000000000000001_0.0001 n2_0.0012000000000000001_0.0001 0
V376 n0_0.0012000000000000001_0.0002 n2_0.0012000000000000001_0.0002 0
V377 n0_0.0012000000000000001_0.00030000000000000003 n2_0.0012000000000000001_0.00030000000000000003 0
V378 n0_0.0012000000000000001_0.0004 n2_0.0012000000000000001_0.0004 0
V379 n0_0.0012000000000000001_0.0005 n2_0.0012000000000000001_0.0005 0
V380 n0_0.0012000000000000001_0.0006000000000000001 n2_0.0012000000000000001_0.0006000000000000001 0
V381 n0_0.0012000000000000001_0.0007 n2_0.0012000000000000001_0.0007 0
V382 n0_0.0012000000000000001_0.0008 n2_0.0012000000000000001_0.0008 0
V383 n0_0.0012000000000000001_0.0009000000000000001 n2_0.0012000000000000001_0.0009000000000000001 0
V384 n0_0.0012000000000000001_0.001 n2_0.0012000000000000001_0.001 0
V385 n0_0.0012000000000000001_0.0011 n2_0.0012000000000000001_0.0011 0
V386 n0_0.0012000000000000001_0.0012000000000000001 n2_0.0012000000000000001_0.0012000000000000001 0
V387 n0_0.0012000000000000001_0.0013000000000000002 n2_0.0012000000000000001_0.0013000000000000002 0
V388 n0_0.0012000000000000001_0.0014 n2_0.0012000000000000001_0.0014 0
V389 n0_0.0012000000000000001_0.0015 n2_0.0012000000000000001_0.0015 0
V390 n0_0.0012000000000000001_0.0016 n2_0.0012000000000000001_0.0016 0
V391 n0_0.0014_0.0 n2_0.0014_0.0 0
V392 n0_0.0014_0.0001 n2_0.0014_0.0001 0
V393 n0_0.0014_0.0002 n2_0.0014_0.0002 0
V394 n0_0.0014_0.00030000000000000003 n2_0.0014_0.00030000000000000003 0
V395 n0_0.0014_0.0004 n2_0.0014_0.0004 0
V396 n0_0.0014_0.0005 n2_0.0014_0.0005 0
V397 n0_0.0014_0.0006000000000000001 n2_0.0014_0.0006000000000000001 0
V398 n0_0.0014_0.0007 n2_0.0014_0.0007 0
V399 n0_0.0014_0.0008 n2_0.0014_0.0008 0
V400 n0_0.0014_0.0009000000000000001 n2_0.0014_0.0009000000000000001 0
V401 n0_0.0014_0.001 n2_0.0014_0.001 0
V402 n0_0.0014_0.0011 n2_0.0014_0.0011 0
V403 n0_0.0014_0.0012000000000000001 n2_0.0014_0.0012000000000000001 0
V404 n0_0.0014_0.0013000000000000002 n2_0.0014_0.0013000000000000002 0
V405 n0_0.0014_0.0014 n2_0.0014_0.0014 0
V406 n0_0.0014_0.0015 n2_0.0014_0.0015 0
V407 n0_0.0014_0.0016 n2_0.0014_0.0016 0
V408 n0_0.0016_0.0 n2_0.0016_0.0 0
V409 n0_0.0016_0.0001 n2_0.0016_0.0001 0
V410 n0_0.0016_0.0002 n2_0.0016_0.0002 0
V411 n0_0.0016_0.00030000000000000003 n2_0.0016_0.00030000000000000003 0
V412 n0_0.0016_0.0004 n2_0.0016_0.0004 0
V413 n0_0.0016_0.0005 n2_0.0016_0.0005 0
V414 n0_0.0016_0.0006000000000000001 n2_0.0016_0.0006000000000000001 0
V415 n0_0.0016_0.0007 n2_0.0016_0.0007 0
V416 n0_0.0016_0.0008 n2_0.0016_0.0008 0
V417 n0_0.0016_0.0009000000000000001 n2_0.0016_0.0009000000000000001 0
V418 n0_0.0016_0.001 n2_0.0016_0.001 0
V419 n0_0.0016_0.0011 n2_0.0016_0.0011 0
V420 n0_0.0016_0.0012000000000000001 n2_0.0016_0.0012000000000000001 0
V421 n0_0.0016_0.0013000000000000002 n2_0.0016_0.0013000000000000002 0
V422 n0_0.0016_0.0014 n2_0.0016_0.0014 0
V423 n0_0.0016_0.0015 n2_0.0016_0.0015 0
V424 n0_0.0016_0.0016 n2_0.0016_0.0016 0
* layer: M2,VDD net: 2
R425 n2_0.0_0.0 n2_0.0_0.0001 0.011008996600000001
R426 n2_0.0_0.0001 n2_0.0_0.0002 0.011008996600000001
R427 n2_0.0_0.0002 n2_0.0_0.00030000000000000003 0.011008996600000001
R428 n2_0.0_0.00030000000000000003 n2_0.0_0.0004 0.011008996600000001
R429 n2_0.0_0.0004 n2_0.0_0.0005 0.011008996600000001
R430 n2_0.0_0.0005 n2_0.0_0.0006000000000000001 0.011008996600000001
R431 n2_0.0_0.0006000000000000001 n2_0.0_0.0007 0.011008996600000001
R432 n2_0.0_0.0007 n2_0.0_0.0008 0.011008996600000001
R433 n2_0.0_0.0008 n2_0.0_0.0009000000000000001 0.011008996600000001
R434 n2_0.0_0.0009000000000000001 n2_0.0_0.001 0.011008996600000001
R435 n2_0.0_0.001 n2_0.0_0.0011 0.011008996600000001
R436 n2_0.0_0.0011 n2_0.0_0.0012000000000000001 0.011008996600000001
R437 n2_0.0_0.0012000000000000001 n2_0.0_0.0013000000000000002 0.011008996600000001
R438 n2_0.0_0.0013000000000000002 n2_0.0_0.0014 0.011008996600000001
R439 n2_0.0_0.0014 n2_0.0_0.0015 0.011008996600000001
R440 n2_0.0_0.0015 n2_0.0_0.0016 0.011008996600000001
R441 n2_0.0002_0.0 n2_0.0002_0.0001 0.011008996600000001
R442 n2_0.0002_0.0001 n2_0.0002_0.0002 0.011008996600000001
R443 n2_0.0002_0.0002 n2_0.0002_0.00030000000000000003 0.011008996600000001
R444 n2_0.0002_0.00030000000000000003 n2_0.0002_0.0004 0.011008996600000001
R445 n2_0.0002_0.0004 n2_0.0002_0.0005 0.011008996600000001
R446 n2_0.0002_0.0005 n2_0.0002_0.0006000000000000001 0.011008996600000001
R447 n2_0.0002_0.0006000000000000001 n2_0.0002_0.0007 0.011008996600000001
R448 n2_0.0002_0.0007 n2_0.0002_0.0008 0.011008996600000001
R449 n2_0.0002_0.0008 n2_0.0002_0.0009000000000000001 0.011008996600000001
R450 n2_0.0002_0.0009000000000000001 n2_0.0002_0.001 0.011008996600000001
R451 n2_0.0002_0.001 n2_0.0002_0.0011 0.011008996600000001
R452 n2_0.0002_0.0011 n2_0.0002_0.0012000000000000001 0.011008996600000001
R453 n2_0.0002_0.0012000000000000001 n2_0.0002_0.0013000000000000002 0.011008996600000001
R454 n2_0.0002_0.0013000000000000002 n2_0.0002_0.0014 0.011008996600000001
R455 n2_0.0002_0.0014 n2_0.0002_0.0015 0.011008996600000001
R456 n2_0.0002_0.0015 n2_0.0002_0.0016 0.011008996600000001
R457 n2_0.0004_0.0 n2_0.0004_0.0001 0.011008996600000001
R458 n2_0.0004_0.0001 n2_0.0004_0.0002 0.011008996600000001
R459 n2_0.0004_0.0002 n2_0.0004_0.00030000000000000003 0.011008996600000001
R460 n2_0.0004_0.00030000000000000003 n2_0.0004_0.0004 0.011008996600000001
R461 n2_0.0004_0.0004 n2_0.0004_0.0005 0.011008996600000001
R462 n2_0.0004_0.0005 n2_0.0004_0.0006000000000000001 0.011008996600000001
R463 n2_0.0004_0.0006000000000000001 n2_0.0004_0.0007 0.011008996600000001
R464 n2_0.0004_0.0007 n2_0.0004_0.0008 0.011008996600000001
R465 n2_0.0004_0.0008 n2_0.0004_0.0009000000000000001 0.011008996600000001
R466 n2_0.0004_0.0009000000000000001 n2_0.0004_0.001 0.011008996600000001
R467 n2_0.0004_0.001 n2_0.0004_0.0011 0.011008996600000001
R468 n2_0.0004_0.0011 n2_0.0004_0.0012000000000000001 0.011008996600000001
R469 n2_0.0004_0.0012000000000000001 n2_0.0004_0.0013000000000000002 0.011008996600000001
R470 n2_0.0004_0.0013000000000000002 n2_0.0004_0.0014 0.011008996600000001
R471 n2_0.0004_0.0014 n2_0.0004_0.0015 0.011008996600000001
R472 n2_0.0004_0.0015 n2_0.0004_0.0016 0.011008996600000001
R473 n2_0.0006000000000000001_0.0 n2_0.0006000000000000001_0.0001 0.011008996600000001
R474 n2_0.0006000000000000001_0.0001 n2_0.0006000000000000001_0.0002 0.011008996600000001
R475 n2_0.0006000000000000001_0.0002 n2_0.0006000000000000001_0.00030000000000000003 0.011008996600000001
R476 n2_0.0006000000000000001_0.00030000000000000003 n2_0.0006000000000000001_0.0004 0.011008996600000001
R477 n2_0.0006000000000000001_0.0004 n2_0.0006000000000000001_0.0005 0.011008996600000001
R478 n2_0.0006000000000000001_0.0005 n2_0.0006000000000000001_0.0006000000000000001 0.011008996600000001
R479 n2_0.0006000000000000001_0.0006000000000000001 n2_0.0006000000000000001_0.0007 0.011008996600000001
R480 n2_0.0006000000000000001_0.0007 n2_0.0006000000000000001_0.0008 0.011008996600000001
R481 n2_0.0006000000000000001_0.0008 n2_0.0006000000000000001_0.0009000000000000001 0.011008996600000001
R482 n2_0.0006000000000000001_0.0009000000000000001 n2_0.0006000000000000001_0.001 0.011008996600000001
R483 n2_0.0006000000000000001_0.001 n2_0.0006000000000000001_0.0011 0.011008996600000001
R484 n2_0.0006000000000000001_0.0011 n2_0.0006000000000000001_0.0012000000000000001 0.011008996600000001
R485 n2_0.0006000000000000001_0.0012000000000000001 n2_0.0006000000000000001_0.0013000000000000002 0.011008996600000001
R486 n2_0.0006000000000000001_0.0013000000000000002 n2_0.0006000000000000001_0.0014 0.011008996600000001
R487 n2_0.0006000000000000001_0.0014 n2_0.0006000000000000001_0.0015 0.011008996600000001
R488 n2_0.0006000000000000001_0.0015 n2_0.0006000000000000001_0.0016 0.011008996600000001
R489 n2_0.0008_0.0 n2_0.0008_0.0001 0.011008996600000001
R490 n2_0.0008_0.0001 n2_0.0008_0.0002 0.011008996600000001
R491 n2_0.0008_0.0002 n2_0.0008_0.00030000000000000003 0.011008996600000001
R492 n2_0.0008_0.00030000000000000003 n2_0.0008_0.0004 0.011008996600000001
R493 n2_0.0008_0.0004 n2_0.0008_0.0005 0.011008996600000001
R494 n2_0.0008_0.0005 n2_0.0008_0.0006000000000000001 0.011008996600000001
R495 n2_0.0008_0.0006000000000000001 n2_0.0008_0.0007 0.011008996600000001
R496 n2_0.0008_0.0007 n2_0.0008_0.0008 0.011008996600000001
R497 n2_0.0008_0.0008 n2_0.0008_0.0009000000000000001 0.011008996600000001
R498 n2_0.0008_0.0009000000000000001 n2_0.0008_0.001 0.011008996600000001
R499 n2_0.0008_0.001 n2_0.0008_0.0011 0.011008996600000001
R500 n2_0.0008_0.0011 n2_0.0008_0.0012000000000000001 0.011008996600000001
R501 n2_0.0008_0.0012000000000000001 n2_0.0008_0.0013000000000000002 0.011008996600000001
R502 n2_0.0008_0.0013000000000000002 n2_0.0008_0.0014 0.011008996600000001
R503 n2_0.0008_0.0014 n2_0.0008_0.0015 0.011008996600000001
R504 n2_0.0008_0.0015 n2_0.0008_0.0016 0.011008996600000001
R505 n2_0.001_0.0 n2_0.001_0.0001 0.011008996600000001
R506 n2_0.001_0.0001 n2_0.001_0.0002 0.011008996600000001
R507 n2_0.001_0.0002 n2_0.001_0.00030000000000000003 0.011008996600000001
R508 n2_0.001_0.00030000000000000003 n2_0.001_0.0004 0.011008996600000001
R509 n2_0.001_0.0004 n2_0.001_0.0005 0.011008996600000001
R510 n2_0.001_0.0005 n2_0.001_0.0006000000000000001 0.011008996600000001
R511 n2_0.001_0.0006000000000000001 n2_0.001_0.0007 0.011008996600000001
R512 n2_0.001_0.0007 n2_0.001_0.0008 0.011008996600000001
R513 n2_0.001_0.0008 n2_0.001_0.0009000000000000001 0.011008996600000001
R514 n2_0.001_0.0009000000000000001 n2_0.001_0.001 0.011008996600000001
R515 n2_0.001_0.001 n2_0.001_0.0011 0.011008996600000001
R516 n2_0.001_0.0011 n2_0.001_0.0012000000000000001 0.011008996600000001
R517 n2_0.001_0.0012000000000000001 n2_0.001_0.0013000000000000002 0.011008996600000001
R518 n2_0.001_0.0013000000000000002 n2_0.001_0.0014 0.011008996600000001
R519 n2_0.001_0.0014 n2_0.001_0.0015 0.011008996600000001
R520 n2_0.001_0.0015 n2_0.001_0.0016 0.011008996600000001
R521 n2_0.0012000000000000001_0.0 n2_0.0012000000000000001_0.0001 0.011008996600000001
R522 n2_0.0012000000000000001_0.0001 n2_0.0012000000000000001_0.0002 0.011008996600000001
R523 n2_0.0012000000000000001_0.0002 n2_0.0012000000000000001_0.00030000000000000003 0.011008996600000001
R524 n2_0.0012000000000000001_0.00030000000000000003 n2_0.0012000000000000001_0.0004 0.011008996600000001
R525 n2_0.0012000000000000001_0.0004 n2_0.0012000000000000001_0.0005 0.011008996600000001
R526 n2_0.0012000000000000001_0.0005 n2_0.0012000000000000001_0.0006000000000000001 0.011008996600000001
R527 n2_0.0012000000000000001_0.0006000000000000001 n2_0.0012000000000000001_0.0007 0.011008996600000001
R528 n2_0.0012000000000000001_0.0007 n2_0.0012000000000000001_0.0008 0.011008996600000001
R529 n2_0.0012000000000000001_0.0008 n2_0.0012000000000000001_0.0009000000000000001 0.011008996600000001
R530 n2_0.0012000000000000001_0.0009000000000000001 n2_0.0012000000000000001_0.001 0.011008996600000001
R531 n2_0.0012000000000000001_0.001 n2_0.0012000000000000001_0.0011 0.011008996600000001
R532 n2_0.0012000000000000001_0.0011 n2_0.0012000000000000001_0.0012000000000000001 0.011008996600000001
R533 n2_0.0012000000000000001_0.0012000000000000001 n2_0.0012000000000000001_0.0013000000000000002 0.011008996600000001
R534 n2_0.0012000000000000001_0.0013000000000000002 n2_0.0012000000000000001_0.0014 0.011008996600000001
R535 n2_0.0012000000000000001_0.0014 n2_0.0012000000000000001_0.0015 0.011008996600000001
R536 n2_0.0012000000000000001_0.0015 n2_0.0012000000000000001_0.0016 0.011008996600000001
R537 n2_0.0014_0.0 n2_0.0014_0.0001 0.011008996600000001
R538 n2_0.0014_0.0001 n2_0.0014_0.0002 0.011008996600000001
R539 n2_0.0014_0.0002 n2_0.0014_0.00030000000000000003 0.011008996600000001
R540 n2_0.0014_0.00030000000000000003 n2_0.0014_0.0004 0.011008996600000001
R541 n2_0.0014_0.0004 n2_0.0014_0.0005 0.011008996600000001
R542 n2_0.0014_0.0005 n2_0.0014_0.0006000000000000001 0.011008996600000001
R543 n2_0.0014_0.0006000000000000001 n2_0.0014_0.0007 0.011008996600000001
R544 n2_0.0014_0.0007 n2_0.0014_0.0008 0.011008996600000001
R545 n2_0.0014_0.0008 n2_0.0014_0.0009000000000000001 0.011008996600000001
R546 n2_0.0014_0.0009000000000000001 n2_0.0014_0.001 0.011008996600000001
R547 n2_0.0014_0.001 n2_0.0014_0.0011 0.011008996600000001
R548 n2_0.0014_0.0011 n2_0.0014_0.0012000000000000001 0.011008996600000001
R549 n2_0.0014_0.0012000000000000001 n2_0.0014_0.0013000000000000002 0.011008996600000001
R550 n2_0.0014_0.0013000000000000002 n2_0.0014_0.0014 0.011008996600000001
R551 n2_0.0014_0.0014 n2_0.0014_0.0015 0.011008996600000001
R552 n2_0.0014_0.0015 n2_0.0014_0.0016 0.011008996600000001
R553 n2_0.0016_0.0 n2_0.0016_0.0001 0.011008996600000001
R554 n2_0.0016_0.0001 n2_0.0016_0.0002 0.011008996600000001
R555 n2_0.0016_0.0002 n2_0.0016_0.00030000000000000003 0.011008996600000001
R556 n2_0.0016_0.00030000000000000003 n2_0.0016_0.0004 0.011008996600000001
R557 n2_0.0016_0.0004 n2_0.0016_0.0005 0.011008996600000001
R558 n2_0.0016_0.0005 n2_0.0016_0.0006000000000000001 0.011008996600000001
R559 n2_0.0016_0.0006000000000000001 n2_0.0016_0.0007 0.011008996600000001
R560 n2_0.0016_0.0007 n2_0.0016_0.0008 0.011008996600000001
R561 n2_0.0016_0.0008 n2_0.0016_0.0009000000000000001 0.011008996600000001
R562 n2_0.0016_0.0009000000000000001 n2_0.0016_0.001 0.011008996600000001
R563 n2_0.0016_0.001 n2_0.0016_0.0011 0.011008996600000001
R564 n2_0.0016_0.0011 n2_0.0016_0.0012000000000000001 0.011008996600000001
R565 n2_0.0016_0.0012000000000000001 n2_0.0016_0.0013000000000000002 0.011008996600000001
R566 n2_0.0016_0.0013000000000000002 n2_0.0016_0.0014 0.011008996600000001
R567 n2_0.0016_0.0014 n2_0.0016_0.0015 0.011008996600000001
R568 n2_0.0016_0.0015 n2_0.0016_0.0016 0.011008996600000001
* vias from: 2 to 4
V569 n2_0.0_0.0 n4_0.0_0.0 0
V570 n2_0.0_0.0002 n4_0.0_0.0002 0
V571 n2_0.0_0.0004 n4_0.0_0.0004 0
V572 n2_0.0_0.0006000000000000001 n4_0.0_0.0006000000000000001 0
V573 n2_0.0_0.0008 n4_0.0_0.0008 0
V574 n2_0.0_0.001 n4_0.0_0.001 0
V575 n2_0.0_0.0012000000000000001 n4_0.0_0.0012000000000000001 0
V576 n2_0.0_0.0014 n4_0.0_0.0014 0
V577 n2_0.0_0.0016 n4_0.0_0.0016 0
V578 n2_0.0002_0.0 n4_0.0002_0.0 0
V579 n2_0.0002_0.0002 n4_0.0002_0.0002 0
V580 n2_0.0002_0.0004 n4_0.0002_0.0004 0
V581 n2_0.0002_0.0006000000000000001 n4_0.0002_0.0006000000000000001 0
V582 n2_0.0002_0.0008 n4_0.0002_0.0008 0
V583 n2_0.0002_0.001 n4_0.0002_0.001 0
V584 n2_0.0002_0.0012000000000000001 n4_0.0002_0.0012000000000000001 0
V585 n2_0.0002_0.0014 n4_0.0002_0.0014 0
V586 n2_0.0002_0.0016 n4_0.0002_0.0016 0
V587 n2_0.0004_0.0 n4_0.0004_0.0 0
V588 n2_0.0004_0.0002 n4_0.0004_0.0002 0
V589 n2_0.0004_0.0004 n4_0.0004_0.0004 0
V590 n2_0.0004_0.0006000000000000001 n4_0.0004_0.0006000000000000001 0
V591 n2_0.0004_0.0008 n4_0.0004_0.0008 0
V592 n2_0.0004_0.001 n4_0.0004_0.001 0
V593 n2_0.0004_0.0012000000000000001 n4_0.0004_0.0012000000000000001 0
V594 n2_0.0004_0.0014 n4_0.0004_0.0014 0
V595 n2_0.0004_0.0016 n4_0.0004_0.0016 0
V596 n2_0.0006000000000000001_0.0 n4_0.0006000000000000001_0.0 0
V597 n2_0.0006000000000000001_0.0002 n4_0.0006000000000000001_0.0002 0
V598 n2_0.0006000000000000001_0.0004 n4_0.0006000000000000001_0.0004 0
V599 n2_0.0006000000000000001_0.0006000000000000001 n4_0.0006000000000000001_0.0006000000000000001 0
V600 n2_0.0006000000000000001_0.0008 n4_0.0006000000000000001_0.0008 0
V601 n2_0.0006000000000000001_0.001 n4_0.0006000000000000001_0.001 0
V602 n2_0.0006000000000000001_0.0012000000000000001 n4_0.0006000000000000001_0.0012000000000000001 0
V603 n2_0.0006000000000000001_0.0014 n4_0.0006000000000000001_0.0014 0
V604 n2_0.0006000000000000001_0.0016 n4_0.0006000000000000001_0.0016 0
V605 n2_0.0008_0.0 n4_0.0008_0.0 0
V606 n2_0.0008_0.0002 n4_0.0008_0.0002 0
V607 n2_0.0008_0.0004 n4_0.0008_0.0004 0
V608 n2_0.0008_0.0006000000000000001 n4_0.0008_0.0006000000000000001 0
V609 n2_0.0008_0.0008 n4_0.0008_0.0008 0
V610 n2_0.0008_0.001 n4_0.0008_0.001 0
V611 n2_0.0008_0.0012000000000000001 n4_0.0008_0.0012000000000000001 0
V612 n2_0.0008_0.0014 n4_0.0008_0.0014 0
V613 n2_0.0008_0.0016 n4_0.0008_0.0016 0
V614 n2_0.001_0.0 n4_0.001_0.0 0
V615 n2_0.001_0.0002 n4_0.001_0.0002 0
V616 n2_0.001_0.0004 n4_0.001_0.0004 0
V617 n2_0.001_0.0006000000000000001 n4_0.001_0.0006000000000000001 0
V618 n2_0.001_0.0008 n4_0.001_0.0008 0
V619 n2_0.001_0.001 n4_0.001_0.001 0
V620 n2_0.001_0.0012000000000000001 n4_0.001_0.0012000000000000001 0
V621 n2_0.001_0.0014 n4_0.001_0.0014 0
V622 n2_0.001_0.0016 n4_0.001_0.0016 0
V623 n2_0.0012000000000000001_0.0 n4_0.0012000000000000001_0.0 0
V624 n2_0.0012000000000000001_0.0002 n4_0.0012000000000000001_0.0002 0
V625 n2_0.0012000000000000001_0.0004 n4_0.0012000000000000001_0.0004 0
V626 n2_0.0012000000000000001_0.0006000000000000001 n4_0.0012000000000000001_0.0006000000000000001 0
V627 n2_0.0012000000000000001_0.0008 n4_0.0012000000000000001_0.0008 0
V628 n2_0.0012000000000000001_0.001 n4_0.0012000000000000001_0.001 0
V629 n2_0.0012000000000000001_0.0012000000000000001 n4_0.0012000000000000001_0.0012000000000000001 0
V630 n2_0.0012000000000000001_0.0014 n4_0.0012000000000000001_0.0014 0
V631 n2_0.0012000000000000001_0.0016 n4_0.0012000000000000001_0.0016 0
V632 n2_0.0014_0.0 n4_0.0014_0.0 0
V633 n2_0.0014_0.0002 n4_0.0014_0.0002 0
V634 n2_0.0014_0.0004 n4_0.0014_0.0004 0
V635 n2_0.0014_0.0006000000000000001 n4_0.0014_0.0006000000000000001 0
V636 n2_0.0014_0.0008 n4_0.0014_0.0008 0
V637 n2_0.0014_0.001 n4_0.0014_0.001 0
V638 n2_0.0014_0.0012000000000000001 n4_0.0014_0.0012000000000000001 0
V639 n2_0.0014_0.0014 n4_0.0014_0.0014 0
V640 n2_0.0014_0.0016 n4_0.0014_0.0016 0
V641 n2_0.0016_0.0 n4_0.0016_0.0 0
V642 n2_0.0016_0.0002 n4_0.0016_0.0002 0
V643 n2_0.0016_0.0004 n4_0.0016_0.0004 0
V644 n2_0.0016_0.0006000000000000001 n4_0.0016_0.0006000000000000001 0
V645 n2_0.0016_0.0008 n4_0.0016_0.0008 0
V646 n2_0.0016_0.001 n4_0.0016_0.001 0
V647 n2_0.0016_0.0012000000000000001 n4_0.0016_0.0012000000000000001 0
V648 n2_0.0016_0.0014 n4_0.0016_0.0014 0
V649 n2_0.0016_0.0016 n4_0.0016_0.0016 0
* layer: M3,VDD net: 4
R650 n4_0.0_0.0 n4_0.0002_0.0 0.019989181600000003
R651 n4_0.0002_0.0 n4_0.0004_0.0 0.019989181600000003
R652 n4_0.0004_0.0 n4_0.0006000000000000001_0.0 0.019989181600000003
R653 n4_0.0006000000000000001_0.0 n4_0.0008_0.0 0.019989181600000003
R654 n4_0.0008_0.0 n4_0.001_0.0 0.019989181600000003
R655 n4_0.001_0.0 n4_0.0012000000000000001_0.0 0.019989181600000003
R656 n4_0.0012000000000000001_0.0 n4_0.0014_0.0 0.019989181600000003
R657 n4_0.0014_0.0 n4_0.0016_0.0 0.019989181600000003
R658 n4_0.0_0.0002 n4_0.0002_0.0002 0.019989181600000003
R659 n4_0.0002_0.0002 n4_0.0004_0.0002 0.019989181600000003
R660 n4_0.0004_0.0002 n4_0.0006000000000000001_0.0002 0.019989181600000003
R661 n4_0.0006000000000000001_0.0002 n4_0.0008_0.0002 0.019989181600000003
R662 n4_0.0008_0.0002 n4_0.001_0.0002 0.019989181600000003
R663 n4_0.001_0.0002 n4_0.0012000000000000001_0.0002 0.019989181600000003
R664 n4_0.0012000000000000001_0.0002 n4_0.0014_0.0002 0.019989181600000003
R665 n4_0.0014_0.0002 n4_0.0016_0.0002 0.019989181600000003
R666 n4_0.0_0.0004 n4_0.0002_0.0004 0.019989181600000003
R667 n4_0.0002_0.0004 n4_0.0004_0.0004 0.019989181600000003
R668 n4_0.0004_0.0004 n4_0.0006000000000000001_0.0004 0.019989181600000003
R669 n4_0.0006000000000000001_0.0004 n4_0.0008_0.0004 0.019989181600000003
R670 n4_0.0008_0.0004 n4_0.001_0.0004 0.019989181600000003
R671 n4_0.001_0.0004 n4_0.0012000000000000001_0.0004 0.019989181600000003
R672 n4_0.0012000000000000001_0.0004 n4_0.0014_0.0004 0.019989181600000003
R673 n4_0.0014_0.0004 n4_0.0016_0.0004 0.019989181600000003
R674 n4_0.0_0.0006000000000000001 n4_0.0002_0.0006000000000000001 0.019989181600000003
R675 n4_0.0002_0.0006000000000000001 n4_0.0004_0.0006000000000000001 0.019989181600000003
R676 n4_0.0004_0.0006000000000000001 n4_0.0006000000000000001_0.0006000000000000001 0.019989181600000003
R677 n4_0.0006000000000000001_0.0006000000000000001 n4_0.0008_0.0006000000000000001 0.019989181600000003
R678 n4_0.0008_0.0006000000000000001 n4_0.001_0.0006000000000000001 0.019989181600000003
R679 n4_0.001_0.0006000000000000001 n4_0.0012000000000000001_0.0006000000000000001 0.019989181600000003
R680 n4_0.0012000000000000001_0.0006000000000000001 n4_0.0014_0.0006000000000000001 0.019989181600000003
R681 n4_0.0014_0.0006000000000000001 n4_0.0016_0.0006000000000000001 0.019989181600000003
R682 n4_0.0_0.0008 n4_0.0002_0.0008 0.019989181600000003
R683 n4_0.0002_0.0008 n4_0.0004_0.0008 0.019989181600000003
R684 n4_0.0004_0.0008 n4_0.0006000000000000001_0.0008 0.019989181600000003
R685 n4_0.0006000000000000001_0.0008 n4_0.0008_0.0008 0.019989181600000003
R686 n4_0.0008_0.0008 n4_0.001_0.0008 0.019989181600000003
R687 n4_0.001_0.0008 n4_0.0012000000000000001_0.0008 0.019989181600000003
R688 n4_0.0012000000000000001_0.0008 n4_0.0014_0.0008 0.019989181600000003
R689 n4_0.0014_0.0008 n4_0.0016_0.0008 0.019989181600000003
R690 n4_0.0_0.001 n4_0.0002_0.001 0.019989181600000003
R691 n4_0.0002_0.001 n4_0.0004_0.001 0.019989181600000003
R692 n4_0.0004_0.001 n4_0.0006000000000000001_0.001 0.019989181600000003
R693 n4_0.0006000000000000001_0.001 n4_0.0008_0.001 0.019989181600000003
R694 n4_0.0008_0.001 n4_0.001_0.001 0.019989181600000003
R695 n4_0.001_0.001 n4_0.0012000000000000001_0.001 0.019989181600000003
R696 n4_0.0012000000000000001_0.001 n4_0.0014_0.001 0.019989181600000003
R697 n4_0.0014_0.001 n4_0.0016_0.001 0.019989181600000003
R698 n4_0.0_0.0012000000000000001 n4_0.0002_0.0012000000000000001 0.019989181600000003
R699 n4_0.0002_0.0012000000000000001 n4_0.0004_0.0012000000000000001 0.019989181600000003
R700 n4_0.0004_0.0012000000000000001 n4_0.0006000000000000001_0.0012000000000000001 0.019989181600000003
R701 n4_0.0006000000000000001_0.0012000000000000001 n4_0.0008_0.0012000000000000001 0.019989181600000003
R702 n4_0.0008_0.0012000000000000001 n4_0.001_0.0012000000000000001 0.019989181600000003
R703 n4_0.001_0.0012000000000000001 n4_0.0012000000000000001_0.0012000000000000001 0.019989181600000003
R704 n4_0.0012000000000000001_0.0012000000000000001 n4_0.0014_0.0012000000000000001 0.019989181600000003
R705 n4_0.0014_0.0012000000000000001 n4_0.0016_0.0012000000000000001 0.019989181600000003
R706 n4_0.0_0.0014 n4_0.0002_0.0014 0.019989181600000003
R707 n4_0.0002_0.0014 n4_0.0004_0.0014 0.019989181600000003
R708 n4_0.0004_0.0014 n4_0.0006000000000000001_0.0014 0.019989181600000003
R709 n4_0.0006000000000000001_0.0014 n4_0.0008_0.0014 0.019989181600000003
R710 n4_0.0008_0.0014 n4_0.001_0.0014 0.019989181600000003
R711 n4_0.001_0.0014 n4_0.0012000000000000001_0.0014 0.019989181600000003
R712 n4_0.0012000000000000001_0.0014 n4_0.0014_0.0014 0.019989181600000003
R713 n4_0.0014_0.0014 n4_0.0016_0.0014 0.019989181600000003
R714 n4_0.0_0.0016 n4_0.0002_0.0016 0.019989181600000003
R715 n4_0.0002_0.0016 n4_0.0004_0.0016 0.019989181600000003
R716 n4_0.0004_0.0016 n4_0.0006000000000000001_0.0016 0.019989181600000003
R717 n4_0.0006000000000000001_0.0016 n4_0.0008_0.0016 0.019989181600000003
R718 n4_0.0008_0.0016 n4_0.001_0.0016 0.019989181600000003
R719 n4_0.001_0.0016 n4_0.0012000000000000001_0.0016 0.019989181600000003
R720 n4_0.0012000000000000001_0.0016 n4_0.0014_0.0016 0.019989181600000003
R721 n4_0.0014_0.0016 n4_0.0016_0.0016 0.019989181600000003
rr722 n4_0.0_0.0 _X_n4_0.0_0.0 0.5
v723 _X_n4_0.0_0.0 0 3.7
rr724 n4_0.0_0.0004 _X_n4_0.0_0.0004 0.5
v725 _X_n4_0.0_0.0004 0 3.7
rr726 n4_0.0_0.0008 _X_n4_0.0_0.0008 0.5
v727 _X_n4_0.0_0.0008 0 3.7
rr728 n4_0.0_0.0012000000000000001 _X_n4_0.0_0.0012000000000000001 0.5
v729 _X_n4_0.0_0.0012000000000000001 0 3.7
rr730 n4_0.0_0.0016 _X_n4_0.0_0.0016 0.5
v731 _X_n4_0.0_0.0016 0 3.7
rr732 n4_0.0004_0.0 _X_n4_0.0004_0.0 0.5
v733 _X_n4_0.0004_0.0 0 3.7
rr734 n4_0.0004_0.0004 _X_n4_0.0004_0.0004 0.5
v735 _X_n4_0.0004_0.0004 0 3.7
rr736 n4_0.0004_0.0008 _X_n4_0.0004_0.0008 0.5
v737 _X_n4_0.0004_0.0008 0 3.7
rr738 n4_0.0004_0.0012000000000000001 _X_n4_0.0004_0.0012000000000000001 0.5
v739 _X_n4_0.0004_0.0012000000000000001 0 3.7
rr740 n4_0.0004_0.0016 _X_n4_0.0004_0.0016 0.5
v741 _X_n4_0.0004_0.0016 0 3.7
rr742 n4_0.0008_0.0 _X_n4_0.0008_0.0 0.5
v743 _X_n4_0.0008_0.0 0 3.7
rr744 n4_0.0008_0.0004 _X_n4_0.0008_0.0004 0.5
v745 _X_n4_0.0008_0.0004 0 3.7
rr746 n4_0.0008_0.0008 _X_n4_0.0008_0.0008 0.5
v747 _X_n4_0.0008_0.0008 0 3.7
rr748 n4_0.0008_0.0012000000000000001 _X_n4_0.0008_0.0012000000000000001 0.5
v749 _X_n4_0.0008_0.0012000000000000001 0 3.7
rr750 n4_0.0008_0.0016 _X_n4_0.0008_0.0016 0.5
v751 _X_n4_0.0008_0.0016 0 3.7
rr752 n4_0.0012000000000000001_0.0 _X_n4_0.0012000000000000001_0.0 0.5
v753 _X_n4_0.0012000000000000001_0.0 0 3.7
rr754 n4_0.0012000000000000001_0.0004 _X_n4_0.0012000000000000001_0.0004 0.5
v755 _X_n4_0.0012000000000000001_0.0004 0 3.7
rr756 n4_0.0012000000000000001_0.0008 _X_n4_0.0012000000000000001_0.0008 0.5
v757 _X_n4_0.0012000000000000001_0.0008 0 3.7
rr758 n4_0.0012000000000000001_0.0012000000000000001 _X_n4_0.0012000000000000001_0.0012000000000000001 0.5
v759 _X_n4_0.0012000000000000001_0.0012000000000000001 0 3.7
rr760 n4_0.0012000000000000001_0.0016 _X_n4_0.0012000000000000001_0.0016 0.5
v761 _X_n4_0.0012000000000000001_0.0016 0 3.7
rr762 n4_0.0016_0.0 _X_n4_0.0016_0.0 0.5
v763 _X_n4_0.0016_0.0 0 3.7
rr764 n4_0.0016_0.0004 _X_n4_0.0016_0.0004 0.5
v765 _X_n4_0.0016_0.0004 0 3.7
rr766 n4_0.0016_0.0008 _X_n4_0.0016_0.0008 0.5
v767 _X_n4_0.0016_0.0008 0 3.7
rr768 n4_0.0016_0.0012000000000000001 _X_n4_0.0016_0.0012000000000000001 0.5
v769 _X_n4_0.0016_0.0012000000000000001 0 3.7
rr770 n4_0.0016_0.0016 _X_n4_0.0016_0.0016 0.5
v771 _X_n4_0.0016_0.0016 0 3.7
iB0_0_v n0_0.0_0.0 0 0.0002788795748083931m
iB0_1_v n0_0.0_0.0001 0 0.0002788795748083931m
iB0_2_v n0_0.0_0.0002 0 0.0006740976315712093m
iB0_3_v n0_0.0_0.00030000000000000003 0 0.0006740976315712093m
iB0_4_v n0_0.0_0.0004 0 0.000148909659548338m
iB0_5_v n0_0.0_0.0005 0 0.000148909659548338m
iB0_6_v n0_0.0_0.0006000000000000001 0 0.0002751733765286159m
iB0_7_v n0_0.0_0.0007 0 0.0002751733765286159m
iB0_8_v n0_0.0_0.0008 0 9.837328401344705e-05m
iB0_9_v n0_0.0_0.0009000000000000001 0 9.837328401344705e-05m
iB0_10_v n0_0.0_0.001 0 0.0005270115425010604m
iB0_11_v n0_0.0_0.0011 0 0.0005270115425010604m
iB0_12_v n0_0.0_0.0012000000000000001 0 0.0004393605877621187m
iB0_13_v n0_0.0_0.0013000000000000002 0 0.0004393605877621187m
iB0_14_v n0_0.0_0.0014 0 0.0009286408256900152m
iB0_15_v n0_0.0_0.0015 0 0.0009286408256900152m
iB0_16_v n0_0.0_0.0016 0 0.0005423980800661486m
iB0_17_v n0_0.0001_0.0 0 0.0002788795748083931m
iB0_18_v n0_0.0001_0.0001 0 0.0002788795748083931m
iB0_19_v n0_0.0001_0.0002 0 0.0006740976315712093m
iB0_20_v n0_0.0001_0.00030000000000000003 0 0.0006740976315712093m
iB0_21_v n0_0.0001_0.0004 0 0.000148909659548338m
iB0_22_v n0_0.0001_0.0005 0 0.000148909659548338m
iB0_23_v n0_0.0001_0.0006000000000000001 0 0.0002751733765286159m
iB0_24_v n0_0.0001_0.0007 0 0.0002751733765286159m
iB0_25_v n0_0.0001_0.0008 0 9.837328401344705e-05m
iB0_26_v n0_0.0001_0.0009000000000000001 0 9.837328401344705e-05m
iB0_27_v n0_0.0001_0.001 0 0.0005270115425010604m
iB0_28_v n0_0.0001_0.0011 0 0.0005270115425010604m
iB0_29_v n0_0.0001_0.0012000000000000001 0 0.0004393605877621187m
iB0_30_v n0_0.0001_0.0013000000000000002 0 0.0004393605877621187m
iB0_31_v n0_0.0001_0.0014 0 0.0009286408256900152m
iB0_32_v n0_0.0001_0.0015 0 0.0009286408256900152m
iB0_33_v n0_0.0001_0.0016 0 0.0005423980800661486m
iB0_34_v n0_0.0002_0.0 0 0.00046279744724569223m
iB0_35_v n0_0.0002_0.0001 0 0.00046279744724569223m
iB0_36_v n0_0.0002_0.0002 0 0.0003370229608410247m
iB0_37_v n0_0.0002_0.00030000000000000003 0 0.0003370229608410247m
iB0_38_v n0_0.0002_0.0004 0 0.0006976089085698285m
iB0_39_v n0_0.0002_0.0005 0 0.0006976089085698285m
iB0_40_v n0_0.0002_0.0006000000000000001 0 0.0003455939440231633m
iB0_41_v n0_0.0002_0.0007 0 0.0003455939440231633m
iB0_42_v n0_0.0002_0.0008 0 0.0007040993640796341m
iB0_43_v n0_0.0002_0.0009000000000000001 0 0.0007040993640796341m
iB0_44_v n0_0.0002_0.001 0 0.00025842991477865323m
iB0_45_v n0_0.0002_0.0011 0 0.00025842991477865323m
iB0_46_v n0_0.0002_0.0012000000000000001 0 0.0002212477583708241m
iB0_47_v n0_0.0002_0.0013000000000000002 0 0.0002212477583708241m
iB0_48_v n0_0.0002_0.0014 0 0.0005870380247032433m
iB0_49_v n0_0.0002_0.0015 0 0.0005870380247032433m
iB0_50_v n0_0.0002_0.0016 0 0.0005423980800661486m
iB0_51_v n0_0.00030000000000000003_0.0 0 0.00046279744724569223m
iB0_52_v n0_0.00030000000000000003_0.0001 0 0.00046279744724569223m
iB0_53_v n0_0.00030000000000000003_0.0002 0 0.0003370229608410247m
iB0_54_v n0_0.00030000000000000003_0.00030000000000000003 0 0.0003370229608410247m
iB0_55_v n0_0.00030000000000000003_0.0004 0 0.0006976089085698285m
iB0_56_v n0_0.00030000000000000003_0.0005 0 0.0006976089085698285m
iB0_57_v n0_0.00030000000000000003_0.0006000000000000001 0 0.0003455939440231633m
iB0_58_v n0_0.00030000000000000003_0.0007 0 0.0003455939440231633m
iB0_59_v n0_0.00030000000000000003_0.0008 0 0.0007040993640796341m
iB0_60_v n0_0.00030000000000000003_0.0009000000000000001 0 0.0007040993640796341m
iB0_61_v n0_0.00030000000000000003_0.001 0 0.00025842991477865323m
iB0_62_v n0_0.00030000000000000003_0.0011 0 0.00025842991477865323m
iB0_63_v n0_0.00030000000000000003_0.0012000000000000001 0 0.0002212477583708241m
iB0_64_v n0_0.00030000000000000003_0.0013000000000000002 0 0.0002212477583708241m
iB0_65_v n0_0.00030000000000000003_0.0014 0 0.0005870380247032433m
iB0_66_v n0_0.00030000000000000003_0.0015 0 0.0005870380247032433m
iB0_67_v n0_0.00030000000000000003_0.0016 0 0.0005423980800661486m
iB0_68_v n0_0.0004_0.0 0 0.0006840636145088835m
iB0_69_v n0_0.0004_0.0001 0 0.0006840636145088835m
iB0_70_v n0_0.0004_0.0002 0 0.00024656237531765605m
iB0_71_v n0_0.0004_0.00030000000000000003 0 0.00024656237531765605m
iB0_72_v n0_0.0004_0.0004 0 0.00041496719366245334m
iB0_73_v n0_0.0004_0.0005 0 0.00041496719366245334m
iB0_74_v n0_0.0004_0.0006000000000000001 0 0.0007030467315758192m
iB0_75_v n0_0.0004_0.0007 0 0.0007030467315758192m
iB0_76_v n0_0.0004_0.0008 0 0.0007919048727834968m
iB0_77_v n0_0.0004_0.0009000000000000001 0 0.0007919048727834968m
iB0_78_v n0_0.0004_0.001 0 0.0009043846340620594m
iB0_79_v n0_0.0004_0.0011 0 0.0009043846340620594m
iB0_80_v n0_0.0004_0.0012000000000000001 0 0.0007629040717803228m
iB0_81_v n0_0.0004_0.0013000000000000002 0 0.0007629040717803228m
iB0_82_v n0_0.0004_0.0014 0 0.00044738458960799665m
iB0_83_v n0_0.0004_0.0015 0 0.00044738458960799665m
iB0_84_v n0_0.0004_0.0016 0 0.0005423980800661486m
iB0_85_v n0_0.0005_0.0 0 0.0006840636145088835m
iB0_86_v n0_0.0005_0.0001 0 0.0006840636145088835m
iB0_87_v n0_0.0005_0.0002 0 0.00024656237531765605m
iB0_88_v n0_0.0005_0.00030000000000000003 0 0.00024656237531765605m
iB0_89_v n0_0.0005_0.0004 0 0.00041496719366245334m
iB0_90_v n0_0.0005_0.0005 0 0.00041496719366245334m
iB0_91_v n0_0.0005_0.0006000000000000001 0 0.0007030467315758192m
iB0_92_v n0_0.0005_0.0007 0 0.0007030467315758192m
iB0_93_v n0_0.0005_0.0008 0 0.0007919048727834968m
iB0_94_v n0_0.0005_0.0009000000000000001 0 0.0007919048727834968m
iB0_95_v n0_0.0005_0.001 0 0.0009043846340620594m
iB0_96_v n0_0.0005_0.0011 0 0.0009043846340620594m
iB0_97_v n0_0.0005_0.0012000000000000001 0 0.0007629040717803228m
iB0_98_v n0_0.0005_0.0013000000000000002 0 0.0007629040717803228m
iB0_99_v n0_0.0005_0.0014 0 0.00044738458960799665m
iB0_100_v n0_0.0005_0.0015 0 0.00044738458960799665m
iB0_101_v n0_0.0005_0.0016 0 0.0005423980800661486m
iB0_102_v n0_0.0006000000000000001_0.0 0 0.0007217064820604806m
iB0_103_v n0_0.0006000000000000001_0.0001 0 0.0007217064820604806m
iB0_104_v n0_0.0006000000000000001_0.0002 0 0.0007521395861772558m
iB0_105_v n0_0.0006000000000000001_0.00030000000000000003 0 0.0007521395861772558m
iB0_106_v n0_0.0006000000000000001_0.0004 0 0.00016855907767689718m
iB0_107_v n0_0.0006000000000000001_0.0005 0 0.00016855907767689718m
iB0_108_v n0_0.0006000000000000001_0.0006000000000000001 0 0.0002939484321308794m
iB0_109_v n0_0.0006000000000000001_0.0007 0 0.0002939484321308794m
iB0_110_v n0_0.0006000000000000001_0.0008 0 0.0005403222905733409m
iB0_111_v n0_0.0006000000000000001_0.0009000000000000001 0 0.0005403222905733409m
iB0_112_v n0_0.0006000000000000001_0.001 0 0.000612340937584976m
iB0_113_v n0_0.0006000000000000001_0.0011 0 0.000612340937584976m
iB0_114_v n0_0.0006000000000000001_0.0012000000000000001 0 0.00045323921772131605m
iB0_115_v n0_0.0006000000000000001_0.0013000000000000002 0 0.00045323921772131605m
iB0_116_v n0_0.0006000000000000001_0.0014 0 0.00023324789719726945m
iB0_117_v n0_0.0006000000000000001_0.0015 0 0.00023324789719726945m
iB0_118_v n0_0.0006000000000000001_0.0016 0 0.0005423980800661486m
iB0_119_v n0_0.0007_0.0 0 0.0007217064820604806m
iB0_120_v n0_0.0007_0.0001 0 0.0007217064820604806m
iB0_121_v n0_0.0007_0.0002 0 0.0007521395861772558m
iB0_122_v n0_0.0007_0.00030000000000000003 0 0.0007521395861772558m
iB0_123_v n0_0.0007_0.0004 0 0.00016855907767689718m
iB0_124_v n0_0.0007_0.0005 0 0.00016855907767689718m
iB0_125_v n0_0.0007_0.0006000000000000001 0 0.0002939484321308794m
iB0_126_v n0_0.0007_0.0007 0 0.0002939484321308794m
iB0_127_v n0_0.0007_0.0008 0 0.0005403222905733409m
iB0_128_v n0_0.0007_0.0009000000000000001 0 0.0005403222905733409m
iB0_129_v n0_0.0007_0.001 0 0.000612340937584976m
iB0_130_v n0_0.0007_0.0011 0 0.000612340937584976m
iB0_131_v n0_0.0007_0.0012000000000000001 0 0.00045323921772131605m
iB0_132_v n0_0.0007_0.0013000000000000002 0 0.00045323921772131605m
iB0_133_v n0_0.0007_0.0014 0 0.00023324789719726945m
iB0_134_v n0_0.0007_0.0015 0 0.00023324789719726945m
iB0_135_v n0_0.0007_0.0016 0 0.0005423980800661486m
iB0_136_v n0_0.0008_0.0 0 0.00035194545467050816m
iB0_137_v n0_0.0008_0.0001 0 0.00035194545467050816m
iB0_138_v n0_0.0008_0.0002 0 0.001000696434567538m
iB0_139_v n0_0.0008_0.00030000000000000003 0 0.001000696434567538m
iB0_140_v n0_0.0008_0.0004 0 0.0004187123012113034m
iB0_141_v n0_0.0008_0.0005 0 0.0004187123012113034m
iB0_142_v n0_0.0008_0.0006000000000000001 0 0.00026906408428224477m
iB0_143_v n0_0.0008_0.0007 0 0.00026906408428224477m
iB0_144_v n0_0.0008_0.0008 0 0.0004255781504248782m
iB0_145_v n0_0.0008_0.0009000000000000001 0 0.0004255781504248782m
iB0_146_v n0_0.0008_0.001 0 0.000554750202491484m
iB0_147_v n0_0.0008_0.0011 0 0.000554750202491484m
iB0_148_v n0_0.0008_0.0012000000000000001 0 0.0006468390661742792m
iB0_149_v n0_0.0008_0.0013000000000000002 0 0.0006468390661742792m
iB0_150_v n0_0.0008_0.0014 0 0.0004570672593667445m
iB0_151_v n0_0.0008_0.0015 0 0.0004570672593667445m
iB0_152_v n0_0.0008_0.0016 0 0.0005423980800661486m
iB0_153_v n0_0.0009000000000000001_0.0 0 0.00035194545467050816m
iB0_154_v n0_0.0009000000000000001_0.0001 0 0.00035194545467050816m
iB0_155_v n0_0.0009000000000000001_0.0002 0 0.001000696434567538m
iB0_156_v n0_0.0009000000000000001_0.00030000000000000003 0 0.001000696434567538m
iB0_157_v n0_0.0009000000000000001_0.0004 0 0.0004187123012113034m
iB0_158_v n0_0.0009000000000000001_0.0005 0 0.0004187123012113034m
iB0_159_v n0_0.0009000000000000001_0.0006000000000000001 0 0.00026906408428224477m
iB0_160_v n0_0.0009000000000000001_0.0007 0 0.00026906408428224477m
iB0_161_v n0_0.0009000000000000001_0.0008 0 0.0004255781504248782m
iB0_162_v n0_0.0009000000000000001_0.0009000000000000001 0 0.0004255781504248782m
iB0_163_v n0_0.0009000000000000001_0.001 0 0.000554750202491484m
iB0_164_v n0_0.0009000000000000001_0.0011 0 0.000554750202491484m
iB0_165_v n0_0.0009000000000000001_0.0012000000000000001 0 0.0006468390661742792m
iB0_166_v n0_0.0009000000000000001_0.0013000000000000002 0 0.0006468390661742792m
iB0_167_v n0_0.0009000000000000001_0.0014 0 0.0004570672593667445m
iB0_168_v n0_0.0009000000000000001_0.0015 0 0.0004570672593667445m
iB0_169_v n0_0.0009000000000000001_0.0016 0 0.0005423980800661486m
iB0_170_v n0_0.001_0.0 0 0.00033606220408432337m
iB0_171_v n0_0.001_0.0001 0 0.00033606220408432337m
iB0_172_v n0_0.001_0.0002 0 0.0005434487807867025m
iB0_173_v n0_0.001_0.00030000000000000003 0 0.0005434487807867025m
iB0_174_v n0_0.001_0.0004 0 0.000665882949620661m
iB0_175_v n0_0.001_0.0005 0 0.000665882949620661m
iB0_176_v n0_0.001_0.0006000000000000001 0 0.000855535523431275m
iB0_177_v n0_0.001_0.0007 0 0.000855535523431275m
iB0_178_v n0_0.001_0.0008 0 0.0003517872379614267m
iB0_179_v n0_0.001_0.0009000000000000001 0 0.0003517872379614267m
iB0_180_v n0_0.001_0.001 0 0.00073919129997313m
iB0_181_v n0_0.001_0.0011 0 0.00073919129997313m
iB0_182_v n0_0.001_0.0012000000000000001 0 0.0002539921783021503m
iB0_183_v n0_0.001_0.0013000000000000002 0 0.0002539921783021503m
iB0_184_v n0_0.001_0.0014 0 0.0004068762273686023m
iB0_185_v n0_0.001_0.0015 0 0.0004068762273686023m
iB0_186_v n0_0.001_0.0016 0 0.0005423980800661486m
iB0_187_v n0_0.0011_0.0 0 0.00033606220408432337m
iB0_188_v n0_0.0011_0.0001 0 0.00033606220408432337m
iB0_189_v n0_0.0011_0.0002 0 0.0005434487807867025m
iB0_190_v n0_0.0011_0.00030000000000000003 0 0.0005434487807867025m
iB0_191_v n0_0.0011_0.0004 0 0.000665882949620661m
iB0_192_v n0_0.0011_0.0005 0 0.000665882949620661m
iB0_193_v n0_0.0011_0.0006000000000000001 0 0.000855535523431275m
iB0_194_v n0_0.0011_0.0007 0 0.000855535523431275m
iB0_195_v n0_0.0011_0.0008 0 0.0003517872379614267m
iB0_196_v n0_0.0011_0.0009000000000000001 0 0.0003517872379614267m
iB0_197_v n0_0.0011_0.001 0 0.00073919129997313m
iB0_198_v n0_0.0011_0.0011 0 0.00073919129997313m
iB0_199_v n0_0.0011_0.0012000000000000001 0 0.0002539921783021503m
iB0_200_v n0_0.0011_0.0013000000000000002 0 0.0002539921783021503m
iB0_201_v n0_0.0011_0.0014 0 0.0004068762273686023m
iB0_202_v n0_0.0011_0.0015 0 0.0004068762273686023m
iB0_203_v n0_0.0011_0.0016 0 0.0005423980800661486m
iB0_204_v n0_0.0012000000000000001_0.0 0 0.00031936961486367426m
iB0_205_v n0_0.0012000000000000001_0.0001 0 0.00031936961486367426m
iB0_206_v n0_0.0012000000000000001_0.0002 0 0.00076521487103465m
iB0_207_v n0_0.0012000000000000001_0.00030000000000000003 0 0.00076521487103465m
iB0_208_v n0_0.0012000000000000001_0.0004 0 0.0007710453577593727m
iB0_209_v n0_0.0012000000000000001_0.0005 0 0.0007710453577593727m
iB0_210_v n0_0.0012000000000000001_0.0006000000000000001 0 0.0004251717796265056m
iB0_211_v n0_0.0012000000000000001_0.0007 0 0.0004251717796265056m
iB0_212_v n0_0.0012000000000000001_0.0008 0 0.0006516894498196907m
iB0_213_v n0_0.0012000000000000001_0.0009000000000000001 0 0.0006516894498196907m
iB0_214_v n0_0.0012000000000000001_0.001 0 0.00012921083715649912m
iB0_215_v n0_0.0012000000000000001_0.0011 0 0.00012921083715649912m
iB0_216_v n0_0.0012000000000000001_0.0012000000000000001 0 0.0002695766312016352m
iB0_217_v n0_0.0012000000000000001_0.0013000000000000002 0 0.0002695766312016352m
iB0_218_v n0_0.0012000000000000001_0.0014 0 0.0008207047082774242m
iB0_219_v n0_0.0012000000000000001_0.0015 0 0.0008207047082774242m
iB0_220_v n0_0.0012000000000000001_0.0016 0 0.0005423980800661486m
iB0_221_v n0_0.0013000000000000002_0.0 0 0.00031936961486367426m
iB0_222_v n0_0.0013000000000000002_0.0001 0 0.00031936961486367426m
iB0_223_v n0_0.0013000000000000002_0.0002 0 0.00076521487103465m
iB0_224_v n0_0.0013000000000000002_0.00030000000000000003 0 0.00076521487103465m
iB0_225_v n0_0.0013000000000000002_0.0004 0 0.0007710453577593727m
iB0_226_v n0_0.0013000000000000002_0.0005 0 0.0007710453577593727m
iB0_227_v n0_0.0013000000000000002_0.0006000000000000001 0 0.0004251717796265056m
iB0_228_v n0_0.0013000000000000002_0.0007 0 0.0004251717796265056m
iB0_229_v n0_0.0013000000000000002_0.0008 0 0.0006516894498196907m
iB0_230_v n0_0.0013000000000000002_0.0009000000000000001 0 0.0006516894498196907m
iB0_231_v n0_0.0013000000000000002_0.001 0 0.00012921083715649912m
iB0_232_v n0_0.0013000000000000002_0.0011 0 0.00012921083715649912m
iB0_233_v n0_0.0013000000000000002_0.0012000000000000001 0 0.0002695766312016352m
iB0_234_v n0_0.0013000000000000002_0.0013000000000000002 0 0.0002695766312016352m
iB0_235_v n0_0.0013000000000000002_0.0014 0 0.0008207047082774242m
iB0_236_v n0_0.0013000000000000002_0.0015 0 0.0008207047082774242m
iB0_237_v n0_0.0013000000000000002_0.0016 0 0.0005423980800661486m
iB0_238_v n0_0.0014_0.0 0 0.0006093219147640054m
iB0_239_v n0_0.0014_0.0001 0 0.0006093219147640054m
iB0_240_v n0_0.0014_0.0002 0 0.0009471622363518463m
iB0_241_v n0_0.0014_0.00030000000000000003 0 0.0009471622363518463m
iB0_242_v n0_0.0014_0.0004 0 0.0003342839631843019m
iB0_243_v n0_0.0014_0.0005 0 0.0003342839631843019m
iB0_244_v n0_0.0014_0.0006000000000000001 0 0.00031724086436300125m
iB0_245_v n0_0.0014_0.0007 0 0.00031724086436300125m
iB0_246_v n0_0.0014_0.0008 0 0.0004660267520651068m
iB0_247_v n0_0.0014_0.0009000000000000001 0 0.0004660267520651068m
iB0_248_v n0_0.0014_0.001 0 2.3362526722990352e-05m
iB0_249_v n0_0.0014_0.0011 0 2.3362526722990352e-05m
iB0_250_v n0_0.0014_0.0012000000000000001 0 3.564358740079494e-05m
iB0_251_v n0_0.0014_0.0013000000000000002 0 3.564358740079494e-05m
iB0_252_v n0_0.0014_0.0014 0 0.0m
iB0_253_v n0_0.0014_0.0015 0 0.0m
iB0_254_v n0_0.0014_0.0016 0 0.0005423980800661486m
iB0_255_v n0_0.0015_0.0 0 0.0006093219147640054m
iB0_256_v n0_0.0015_0.0001 0 0.0006093219147640054m
iB0_257_v n0_0.0015_0.0002 0 0.0009471622363518463m
iB0_258_v n0_0.0015_0.00030000000000000003 0 0.0009471622363518463m
iB0_259_v n0_0.0015_0.0004 0 0.0003342839631843019m
iB0_260_v n0_0.0015_0.0005 0 0.0003342839631843019m
iB0_261_v n0_0.0015_0.0006000000000000001 0 0.00031724086436300125m
iB0_262_v n0_0.0015_0.0007 0 0.00031724086436300125m
iB0_263_v n0_0.0015_0.0008 0 0.0004660267520651068m
iB0_264_v n0_0.0015_0.0009000000000000001 0 0.0004660267520651068m
iB0_265_v n0_0.0015_0.001 0 2.3362526722990352e-05m
iB0_266_v n0_0.0015_0.0011 0 2.3362526722990352e-05m
iB0_267_v n0_0.0015_0.0012000000000000001 0 3.564358740079494e-05m
iB0_268_v n0_0.0015_0.0013000000000000002 0 3.564358740079494e-05m
iB0_269_v n0_0.0015_0.0014 0 0.0m
iB0_270_v n0_0.0015_0.0015 0 0.0m
iB0_271_v n0_0.0015_0.0016 0 0.0005423980800661486m
iB0_272_v n0_0.0016_0.0 0 0.0005423980800661486m
iB0_273_v n0_0.0016_0.0001 0 0.0005423980800661486m
iB0_274_v n0_0.0016_0.0002 0 0.0005423980800661486m
iB0_275_v n0_0.0016_0.00030000000000000003 0 0.0005423980800661486m
iB0_276_v n0_0.0016_0.0004 0 0.0005423980800661486m
iB0_277_v n0_0.0016_0.0005 0 0.0005423980800661486m
iB0_278_v n0_0.0016_0.0006000000000000001 0 0.0005423980800661486m
iB0_279_v n0_0.0016_0.0007 0 0.0005423980800661486m
iB0_280_v n0_0.0016_0.0008 0 0.0005423980800661486m
iB0_281_v n0_0.0016_0.0009000000000000001 0 0.0005423980800661486m
iB0_282_v n0_0.0016_0.001 0 0.0005423980800661486m
iB0_283_v n0_0.0016_0.0011 0 0.0005423980800661486m
iB0_284_v n0_0.0016_0.0012000000000000001 0 0.0005423980800661486m
iB0_285_v n0_0.0016_0.0013000000000000002 0 0.0005423980800661486m
iB0_286_v n0_0.0016_0.0014 0 0.0005423980800661486m
iB0_287_v n0_0.0016_0.0015 0 0.0005423980800661486m
iB0_288_v n0_0.0016_0.0016 0 0.0005423980800661486m
.op
.end